../../../TheSDK_generators/verilog/tb_halfband.v