../../../TheSDK_generators/verilog/halfband.v